TP #3
