TP #1
