TP #2
